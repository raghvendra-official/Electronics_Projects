** Profile: "SCHEMATIC1-SISO"  [ c:\users\raghv\onedrive\desktop\vivado\design1-pspicefiles\schematic1\siso.sim ] 

** Creating circuit file "SISO.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\raghv\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/23.1.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20us 0 
.OPTIONS ADVCONV
.OPTIONS DIGINITSTATE= 0
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
